module ScanCodeToASCII(
    input [7:0] scan_code,
    output [7:0] ascii_code
);
// a	0x61	0x1C	0xF0 0x1C
// b	0x62	0x32	0xF0 0x32
// c	0x63	0x21	0xF0 0x21
// d	0x64	0x23	0xF0 0x23
// e	0x65	0x24	0xF0 0x24
// f	0x66	0x2B	0xF0 0x2B
// g	0x67	0x34	0xF0 0x34
// h	0x68	0x33	0xF0 0x33
// i	0x69	0x43	0xF0 0x43
// j	0x6A	0x3B	0xF0 0x3B
// k	0x6B	0x42	0xF0 0x42
// l	0x6C	0x4B	0xF0 0x4B
// m	0x6D	0x3A	0xF0 0x3A
// n	0x6E	0x31	0xF0 0x31
// o	0x6F	0x44	0xF0 0x44
// p	0x70	0x4D	0xF0 0x4D
// q	0x71	0x15	0xF0 0x15
// r	0x72	0x2D	0xF0 0x2D
// s	0x73	0x1B	0xF0 0x1B
// t	0x74	0x2C	0xF0 0x2C
// u	0x75	0x3C	0xF0 0x3C
// v	0x76	0x2A	0xF0 0x2A
// w	0x77	0x1D	0xF0 0x1D
// x	0x78	0x22	0xF0 0x22
// y	0x79	0x35	0xF0 0x35
// z	0x7A	0x1A	0xF0 0x1A
    MuxKeyWithDefault #(26, 8, 8) ins(
        .out(ascii_code),
        .key(scan_code),
        .default_out(8'hFF),
        .lut({
            8'h1c, 8'h61,
            8'h32, 8'h62,
            8'h21, 8'h63,
            8'h23, 8'h64,
            8'h24, 8'h65,
            8'h2b, 8'h66,
            8'h34, 8'h67,
            8'h33, 8'h68,
            8'h43, 8'h69,
            8'h3b, 8'h6a,
            8'h42, 8'h6b,
            8'h4b, 8'h6c,
            8'h3a, 8'h6d,
            8'h31, 8'h6e,
            8'h44, 8'h6f,
            8'h4d, 8'h70,
            8'h15, 8'h71,
            8'h2d, 8'h72,
            8'h1b, 8'h73,
            8'h2c, 8'h74,
            8'h3c, 8'h75,
            8'h2a, 8'h76,
            8'h1d, 8'h77,
            8'h22, 8'h78,
            8'h35, 8'h79,
            8'h1a, 8'h7a
        })
    );

endmodule //ScanCodeToASCII

